package instNamePackage is
	type instruction_TYPE is (R_ADD, I_ADDI, I_ADDIU, R_ADDU, R_AND, I_ANDI, I_BEQ, I_BNE, J_J ,J_JAL, R_JR, I_LBU, I_LHU, 
		I_LUI, I_LW, NOP, R_NOR, R_OR, I_ORI, R_SLT, I_SLTI, I_SLTIU, R_SLTU, R_SLL, R_SRL, I_SB, I_SH, I_SW, R_SUB, R_SUBU
	);
end instNamePackage;

package body instNamePackage is
	
end instNamePackage;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity hazardUnit is
	port (
		clk : in std_logic;
		rst : in std_logic
	);
end entity hazardUnit;

architecture RTL of hazardUnit is
	
begin

end architecture RTL;
